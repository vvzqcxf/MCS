
.title Vvoltage mode Sensing amplifier 
*****************************
**     Library setting     **
*****************************
.protect
.include '7nm_TT.pm'
.unprotect 

*****************************
**   Circuit Description   **
*****************************
*** By default, m = 1 ***
*** for 1:1:1, the "m" of mos must equal to 1 ***


.subckt SRAM q  qb WL	BL  BLB    

Mpr  q   qb  VDD  x  pmos_sram  m=100
Mnr  q   qb  GND  x  nmos_sram  m=100

Mpl  qb  q  VDD  x  pmos_sram  m=100
Mnl  qb  q  GND  x  nmos_sram  m=100

Mnpr BL  WL  q    x  nmos_sram  m=200
Mnpl BLB WL  qb   x  nmos_sram  m=200

.ends

*****************************
****Precharge Circuit Description***
*****************************

Mp_prel BL    pre   vdd x pmos_sram m=6000
Mp_prer BLB  pre   vdd x pmos_sram m=6000
Mp_pre  BLB  BL pre x pmos_sram m=6000


*****************************
****SA Circuit Description***
*****************************
x1	q0	qb WL_ON	BL	BLB	SRAM

Mpl_top sense    SA_EN     BL     x pmos_sram m=1000
Mpr_top sense_b  SA_EN     BLB    x pmos_sram m=1000
Mpl_mid sense_b  sense     vdd    x pmos_sram m=1000
Mpr_mid sense    sense_b   vdd    x pmos_sram m=1000
Mnl_mid sense_b  sense     mid    x nmos_sram m=2000
Mnr_mid sense    sense_b   mid    x nmos_sram m=2000
Mn_out  mid      SA_EN     gnd    x nmos_sram m=2000



*Mp_pre1l sense    pre   vdd x pmos_sram m=1000
*Mp_pre1r sense_b  pre   vdd x pmos_sram m=1000
*Mp_pr1e  sense_b  sense pre x pmos_sram m=1000


*****************************
**     Voltage Source      **
*****************************
.global VDD GND
.PARAM  BITCAP=1E-12

VVDD VDD GND 0.7v

CBLB BLB GND 512p
CBL  BL  GND 512p

.ic V(BL) =0.7V  
.ic V(BLB)=0.7V  
.ic	V(q0)=0v


VWL_on  WL_on  GND PULSE  ( 0V  0.7V  3ns  0.05ns  0.05ns  0.5ns  1ns )
Vpre  pre  GND PULSE  ( 0V  0.7V  3ns  0.05ns  0.05ns  0.6ns  1ns )
VSAE   SA_EN    GND PULSE  ( 0V  0.7V  3.45ns  0.05ns  0.05ns  0.1ns  1ns )

*****************************
**    Simulator setting    **
*****************************
***************************************
**              option ctrl          **
***************************************
.op
.option post 
.options probe
.probe v(*) i(*)
.tran 0.05ns 25ns

.measure tp_senseEnabletoSense
+ TRIG v(SA_EN) VAL='0.35' RISE=1
+ TARG v(sense) VAL='0.35' fall=1

.measure TRAN Avg_read_pwr  avg POWER from= 3n to=25n




.end


///////////////////////////////////////////////////
.title VM SA 
*****************************
**     Library setting     **
*****************************
.protect
.include '7nm_TT.pm'
.unprotect 
*****************************
**   Circuit Description   **
*****************************
Mpre0 BL  PRE VDD VDD pmos_rvt m=1
Mpre1 BLB PRE VDD VDD pmos_rvt m=1
Mpre2 BL  PRE BLB VDD pmos_rvt m=1
//SRAM
    X0 VDD GND WL[0] BL BLB SRAM        
    X1 VDD GND WL[1] BL BLB SRAM
    X2 VDD GND WL[2] BL BLB SRAM
    X3 VDD GND WL[3] BL BLB SRAM
    X4 VDD GND WL[4] BL BLB SRAM
    X5 VDD GND WL[5] BL BLB SRAM
    X6 VDD GND WL[6] BL BLB SRAM
    X7 VDD GND WL[7] BL BLB SRAM
    X8 VDD GND WL[8] BL BLB SRAM
    X9 VDD GND WL[9] BL BLB SRAM
    X10 VDD GND WL[10] BL BLB SRAM
    X11 VDD GND WL[11] BL BLB SRAM
    X12 VDD GND WL[12] BL BLB SRAM
    X13 VDD GND WL[13] BL BLB SRAM
    X14 VDD GND WL[14] BL BLB SRAM
    X15 VDD GND WL[15] BL BLB SRAM
    X16 VDD GND WL[16] BL BLB SRAM
    X17 VDD GND WL[17] BL BLB SRAM
    X18 VDD GND WL[18] BL BLB SRAM
    X19 VDD GND WL[19] BL BLB SRAM
    X20 VDD GND WL[20] BL BLB SRAM
    X21 VDD GND WL[21] BL BLB SRAM
    X22 VDD GND WL[22] BL BLB SRAM
    X23 VDD GND WL[23] BL BLB SRAM
    X24 VDD GND WL[24] BL BLB SRAM
    X25 VDD GND WL[25] BL BLB SRAM
    X26 VDD GND WL[26] BL BLB SRAM
    X27 VDD GND WL[27] BL BLB SRAM
    X28 VDD GND WL[28] BL BLB SRAM
    X29 VDD GND WL[29] BL BLB SRAM
    X30 VDD GND WL[30] BL BLB SRAM
    X31 VDD GND WL[31] BL BLB SRAM
    X32 VDD GND WL[32] BL BLB SRAM
    X33 VDD GND WL[33] BL BLB SRAM
    X34 VDD GND WL[34] BL BLB SRAM
    X35 VDD GND WL[35] BL BLB SRAM
    X36 VDD GND WL[36] BL BLB SRAM
    X37 VDD GND WL[37] BL BLB SRAM
    X38 VDD GND WL[38] BL BLB SRAM
    X39 VDD GND WL[39] BL BLB SRAM
    X40 VDD GND WL[40] BL BLB SRAM
    X41 VDD GND WL[41] BL BLB SRAM
    X42 VDD GND WL[42] BL BLB SRAM
    X43 VDD GND WL[43] BL BLB SRAM
    X44 VDD GND WL[44] BL BLB SRAM
    X45 VDD GND WL[45] BL BLB SRAM
    X46 VDD GND WL[46] BL BLB SRAM
    X47 VDD GND WL[47] BL BLB SRAM
    X48 VDD GND WL[48] BL BLB SRAM
    X49 VDD GND WL[49] BL BLB SRAM
    X50 VDD GND WL[50] BL BLB SRAM
    X51 VDD GND WL[51] BL BLB SRAM
    X52 VDD GND WL[52] BL BLB SRAM
    X53 VDD GND WL[53] BL BLB SRAM
    X54 VDD GND WL[54] BL BLB SRAM
    X55 VDD GND WL[55] BL BLB SRAM
    X56 VDD GND WL[56] BL BLB SRAM
    X57 VDD GND WL[57] BL BLB SRAM
    X58 VDD GND WL[58] BL BLB SRAM
    X59 VDD GND WL[59] BL BLB SRAM
    X60 VDD GND WL[60] BL BLB SRAM
    X61 VDD GND WL[61] BL BLB SRAM
    X62 VDD GND WL[62] BL BLB SRAM
    X63 VDD GND WL[63] BL BLB SRAM
    X64 VDD GND WL[64] BL BLB SRAM
    X65 VDD GND WL[65] BL BLB SRAM
    X66 VDD GND WL[66] BL BLB SRAM
    X67 VDD GND WL[67] BL BLB SRAM
    X68 VDD GND WL[68] BL BLB SRAM
    X69 VDD GND WL[69] BL BLB SRAM
    X70 VDD GND WL[70] BL BLB SRAM
    X71 VDD GND WL[71] BL BLB SRAM
    X72 VDD GND WL[72] BL BLB SRAM
    X73 VDD GND WL[73] BL BLB SRAM
    X74 VDD GND WL[74] BL BLB SRAM
    X75 VDD GND WL[75] BL BLB SRAM
    X76 VDD GND WL[76] BL BLB SRAM
    X77 VDD GND WL[77] BL BLB SRAM
    X78 VDD GND WL[78] BL BLB SRAM
    X79 VDD GND WL[79] BL BLB SRAM
    X80 VDD GND WL[80] BL BLB SRAM
    X81 VDD GND WL[81] BL BLB SRAM
    X82 VDD GND WL[82] BL BLB SRAM
    X83 VDD GND WL[83] BL BLB SRAM
    X84 VDD GND WL[84] BL BLB SRAM
    X85 VDD GND WL[85] BL BLB SRAM
    X86 VDD GND WL[86] BL BLB SRAM
    X87 VDD GND WL[87] BL BLB SRAM
    X88 VDD GND WL[88] BL BLB SRAM
    X89 VDD GND WL[89] BL BLB SRAM
    X90 VDD GND WL[90] BL BLB SRAM
    X91 VDD GND WL[91] BL BLB SRAM
    X92 VDD GND WL[92] BL BLB SRAM
    X93 VDD GND WL[93] BL BLB SRAM
    X94 VDD GND WL[94] BL BLB SRAM
    X95 VDD GND WL[95] BL BLB SRAM
    X96 VDD GND WL[96] BL BLB SRAM
    X97 VDD GND WL[97] BL BLB SRAM
    X98 VDD GND WL[98] BL BLB SRAM
    X99 VDD GND WL[99] BL BLB SRAM
    X100 VDD GND WL[100] BL BLB SRAM
    X101 VDD GND WL[101] BL BLB SRAM
    X102 VDD GND WL[102] BL BLB SRAM
    X103 VDD GND WL[103] BL BLB SRAM
    X104 VDD GND WL[104] BL BLB SRAM
    X105 VDD GND WL[105] BL BLB SRAM
    X106 VDD GND WL[106] BL BLB SRAM
    X107 VDD GND WL[107] BL BLB SRAM
    X108 VDD GND WL[108] BL BLB SRAM
    X109 VDD GND WL[109] BL BLB SRAM
    X110 VDD GND WL[110] BL BLB SRAM
    X111 VDD GND WL[111] BL BLB SRAM
    X112 VDD GND WL[112] BL BLB SRAM
    X113 VDD GND WL[113] BL BLB SRAM
    X114 VDD GND WL[114] BL BLB SRAM
    X115 VDD GND WL[115] BL BLB SRAM
    X116 VDD GND WL[116] BL BLB SRAM
    X117 VDD GND WL[117] BL BLB SRAM
    X118 VDD GND WL[118] BL BLB SRAM
    X119 VDD GND WL[119] BL BLB SRAM
    X120 VDD GND WL[120] BL BLB SRAM
    X121 VDD GND WL[121] BL BLB SRAM
    X122 VDD GND WL[122] BL BLB SRAM
    X123 VDD GND WL[123] BL BLB SRAM
    X124 VDD GND WL[124] BL BLB SRAM
    X125 VDD GND WL[125] BL BLB SRAM
    X126 VDD GND WL[126] BL BLB SRAM
    X127 VDD GND WL[127] BL BLB SRAM
    X128 VDD GND WL[128] BL BLB SRAM
    X129 VDD GND WL[129] BL BLB SRAM
    X130 VDD GND WL[130] BL BLB SRAM
    X131 VDD GND WL[131] BL BLB SRAM
    X132 VDD GND WL[132] BL BLB SRAM
    X133 VDD GND WL[133] BL BLB SRAM
    X134 VDD GND WL[134] BL BLB SRAM
    X135 VDD GND WL[135] BL BLB SRAM
    X136 VDD GND WL[136] BL BLB SRAM
    X137 VDD GND WL[137] BL BLB SRAM
    X138 VDD GND WL[138] BL BLB SRAM
    X139 VDD GND WL[139] BL BLB SRAM
    X140 VDD GND WL[140] BL BLB SRAM
    X141 VDD GND WL[141] BL BLB SRAM
    X142 VDD GND WL[142] BL BLB SRAM
    X143 VDD GND WL[143] BL BLB SRAM
    X144 VDD GND WL[144] BL BLB SRAM
    X145 VDD GND WL[145] BL BLB SRAM
    X146 VDD GND WL[146] BL BLB SRAM
    X147 VDD GND WL[147] BL BLB SRAM
    X148 VDD GND WL[148] BL BLB SRAM
    X149 VDD GND WL[149] BL BLB SRAM
    X150 VDD GND WL[150] BL BLB SRAM
    X151 VDD GND WL[151] BL BLB SRAM
    X152 VDD GND WL[152] BL BLB SRAM
    X153 VDD GND WL[153] BL BLB SRAM
    X154 VDD GND WL[154] BL BLB SRAM
    X155 VDD GND WL[155] BL BLB SRAM
    X156 VDD GND WL[156] BL BLB SRAM
    X157 VDD GND WL[157] BL BLB SRAM
    X158 VDD GND WL[158] BL BLB SRAM
    X159 VDD GND WL[159] BL BLB SRAM
    X160 VDD GND WL[160] BL BLB SRAM
    X161 VDD GND WL[161] BL BLB SRAM
    X162 VDD GND WL[162] BL BLB SRAM
    X163 VDD GND WL[163] BL BLB SRAM
    X164 VDD GND WL[164] BL BLB SRAM
    X165 VDD GND WL[165] BL BLB SRAM
    X166 VDD GND WL[166] BL BLB SRAM
    X167 VDD GND WL[167] BL BLB SRAM
    X168 VDD GND WL[168] BL BLB SRAM
    X169 VDD GND WL[169] BL BLB SRAM
    X170 VDD GND WL[170] BL BLB SRAM
    X171 VDD GND WL[171] BL BLB SRAM
    X172 VDD GND WL[172] BL BLB SRAM
    X173 VDD GND WL[173] BL BLB SRAM
    X174 VDD GND WL[174] BL BLB SRAM
    X175 VDD GND WL[175] BL BLB SRAM
    X176 VDD GND WL[176] BL BLB SRAM
    X177 VDD GND WL[177] BL BLB SRAM
    X178 VDD GND WL[178] BL BLB SRAM
    X179 VDD GND WL[179] BL BLB SRAM
    X180 VDD GND WL[180] BL BLB SRAM
    X181 VDD GND WL[181] BL BLB SRAM
    X182 VDD GND WL[182] BL BLB SRAM
    X183 VDD GND WL[183] BL BLB SRAM
    X184 VDD GND WL[184] BL BLB SRAM
    X185 VDD GND WL[185] BL BLB SRAM
    X186 VDD GND WL[186] BL BLB SRAM
    X187 VDD GND WL[187] BL BLB SRAM
    X188 VDD GND WL[188] BL BLB SRAM
    X189 VDD GND WL[189] BL BLB SRAM
    X190 VDD GND WL[190] BL BLB SRAM
    X191 VDD GND WL[191] BL BLB SRAM
    X192 VDD GND WL[192] BL BLB SRAM
    X193 VDD GND WL[193] BL BLB SRAM
    X194 VDD GND WL[194] BL BLB SRAM
    X195 VDD GND WL[195] BL BLB SRAM
    X196 VDD GND WL[196] BL BLB SRAM
    X197 VDD GND WL[197] BL BLB SRAM
    X198 VDD GND WL[198] BL BLB SRAM
    X199 VDD GND WL[199] BL BLB SRAM
    X200 VDD GND WL[200] BL BLB SRAM
    X201 VDD GND WL[201] BL BLB SRAM
    X202 VDD GND WL[202] BL BLB SRAM
    X203 VDD GND WL[203] BL BLB SRAM
    X204 VDD GND WL[204] BL BLB SRAM
    X205 VDD GND WL[205] BL BLB SRAM
    X206 VDD GND WL[206] BL BLB SRAM
    X207 VDD GND WL[207] BL BLB SRAM
    X208 VDD GND WL[208] BL BLB SRAM
    X209 VDD GND WL[209] BL BLB SRAM
    X210 VDD GND WL[210] BL BLB SRAM
    X211 VDD GND WL[211] BL BLB SRAM
    X212 VDD GND WL[212] BL BLB SRAM
    X213 VDD GND WL[213] BL BLB SRAM
    X214 VDD GND WL[214] BL BLB SRAM
    X215 VDD GND WL[215] BL BLB SRAM
    X216 VDD GND WL[216] BL BLB SRAM
    X217 VDD GND WL[217] BL BLB SRAM
    X218 VDD GND WL[218] BL BLB SRAM
    X219 VDD GND WL[219] BL BLB SRAM
    X220 VDD GND WL[220] BL BLB SRAM
    X221 VDD GND WL[221] BL BLB SRAM
    X222 VDD GND WL[222] BL BLB SRAM
    X223 VDD GND WL[223] BL BLB SRAM
    X224 VDD GND WL[224] BL BLB SRAM
    X225 VDD GND WL[225] BL BLB SRAM
    X226 VDD GND WL[226] BL BLB SRAM
    X227 VDD GND WL[227] BL BLB SRAM
    X228 VDD GND WL[228] BL BLB SRAM
    X229 VDD GND WL[229] BL BLB SRAM
    X230 VDD GND WL[230] BL BLB SRAM
    X231 VDD GND WL[231] BL BLB SRAM
    X232 VDD GND WL[232] BL BLB SRAM
    X233 VDD GND WL[233] BL BLB SRAM
    X234 VDD GND WL[234] BL BLB SRAM
    X235 VDD GND WL[235] BL BLB SRAM
    X236 VDD GND WL[236] BL BLB SRAM
    X237 VDD GND WL[237] BL BLB SRAM
    X238 VDD GND WL[238] BL BLB SRAM
    X239 VDD GND WL[239] BL BLB SRAM
    X240 VDD GND WL[240] BL BLB SRAM
    X241 VDD GND WL[241] BL BLB SRAM
    X242 VDD GND WL[242] BL BLB SRAM
    X243 VDD GND WL[243] BL BLB SRAM
    X244 VDD GND WL[244] BL BLB SRAM
    X245 VDD GND WL[245] BL BLB SRAM
    X246 VDD GND WL[246] BL BLB SRAM
    X247 VDD GND WL[247] BL BLB SRAM
    X248 VDD GND WL[248] BL BLB SRAM
    X249 VDD GND WL[249] BL BLB SRAM
    X250 VDD GND WL[250] BL BLB SRAM
    X251 VDD GND WL[251] BL BLB SRAM
    X252 VDD GND WL[252] BL BLB SRAM
    X253 VDD GND WL[253] BL BLB SRAM
    X254 VDD GND WL[254] BL BLB SRAM
    X255 VDD GND WL[255] BL BLB SRAM
    X256 VDD GND WL[256] BL BLB SRAM
    X257 VDD GND WL[257] BL BLB SRAM
    X258 VDD GND WL[258] BL BLB SRAM
    X259 VDD GND WL[259] BL BLB SRAM
    X260 VDD GND WL[260] BL BLB SRAM
    X261 VDD GND WL[261] BL BLB SRAM
    X262 VDD GND WL[262] BL BLB SRAM
    X263 VDD GND WL[263] BL BLB SRAM
    X264 VDD GND WL[264] BL BLB SRAM
    X265 VDD GND WL[265] BL BLB SRAM
    X266 VDD GND WL[266] BL BLB SRAM
    X267 VDD GND WL[267] BL BLB SRAM
    X268 VDD GND WL[268] BL BLB SRAM
    X269 VDD GND WL[269] BL BLB SRAM
    X270 VDD GND WL[270] BL BLB SRAM
    X271 VDD GND WL[271] BL BLB SRAM
    X272 VDD GND WL[272] BL BLB SRAM
    X273 VDD GND WL[273] BL BLB SRAM
    X274 VDD GND WL[274] BL BLB SRAM
    X275 VDD GND WL[275] BL BLB SRAM
    X276 VDD GND WL[276] BL BLB SRAM
    X277 VDD GND WL[277] BL BLB SRAM
    X278 VDD GND WL[278] BL BLB SRAM
    X279 VDD GND WL[279] BL BLB SRAM
    X280 VDD GND WL[280] BL BLB SRAM
    X281 VDD GND WL[281] BL BLB SRAM
    X282 VDD GND WL[282] BL BLB SRAM
    X283 VDD GND WL[283] BL BLB SRAM
    X284 VDD GND WL[284] BL BLB SRAM
    X285 VDD GND WL[285] BL BLB SRAM
    X286 VDD GND WL[286] BL BLB SRAM
    X287 VDD GND WL[287] BL BLB SRAM
    X288 VDD GND WL[288] BL BLB SRAM
    X289 VDD GND WL[289] BL BLB SRAM
    X290 VDD GND WL[290] BL BLB SRAM
    X291 VDD GND WL[291] BL BLB SRAM
    X292 VDD GND WL[292] BL BLB SRAM
    X293 VDD GND WL[293] BL BLB SRAM
    X294 VDD GND WL[294] BL BLB SRAM
    X295 VDD GND WL[295] BL BLB SRAM
    X296 VDD GND WL[296] BL BLB SRAM
    X297 VDD GND WL[297] BL BLB SRAM
    X298 VDD GND WL[298] BL BLB SRAM
    X299 VDD GND WL[299] BL BLB SRAM
    X300 VDD GND WL[300] BL BLB SRAM
    X301 VDD GND WL[301] BL BLB SRAM
    X302 VDD GND WL[302] BL BLB SRAM
    X303 VDD GND WL[303] BL BLB SRAM
    X304 VDD GND WL[304] BL BLB SRAM
    X305 VDD GND WL[305] BL BLB SRAM
    X306 VDD GND WL[306] BL BLB SRAM
    X307 VDD GND WL[307] BL BLB SRAM
    X308 VDD GND WL[308] BL BLB SRAM
    X309 VDD GND WL[309] BL BLB SRAM
    X310 VDD GND WL[310] BL BLB SRAM
    X311 VDD GND WL[311] BL BLB SRAM
    X312 VDD GND WL[312] BL BLB SRAM
    X313 VDD GND WL[313] BL BLB SRAM
    X314 VDD GND WL[314] BL BLB SRAM
    X315 VDD GND WL[315] BL BLB SRAM
    X316 VDD GND WL[316] BL BLB SRAM
    X317 VDD GND WL[317] BL BLB SRAM
    X318 VDD GND WL[318] BL BLB SRAM
    X319 VDD GND WL[319] BL BLB SRAM
    X320 VDD GND WL[320] BL BLB SRAM
    X321 VDD GND WL[321] BL BLB SRAM
    X322 VDD GND WL[322] BL BLB SRAM
    X323 VDD GND WL[323] BL BLB SRAM
    X324 VDD GND WL[324] BL BLB SRAM
    X325 VDD GND WL[325] BL BLB SRAM
    X326 VDD GND WL[326] BL BLB SRAM
    X327 VDD GND WL[327] BL BLB SRAM
    X328 VDD GND WL[328] BL BLB SRAM
    X329 VDD GND WL[329] BL BLB SRAM
    X330 VDD GND WL[330] BL BLB SRAM
    X331 VDD GND WL[331] BL BLB SRAM
    X332 VDD GND WL[332] BL BLB SRAM
    X333 VDD GND WL[333] BL BLB SRAM
    X334 VDD GND WL[334] BL BLB SRAM
    X335 VDD GND WL[335] BL BLB SRAM
    X336 VDD GND WL[336] BL BLB SRAM
    X337 VDD GND WL[337] BL BLB SRAM
    X338 VDD GND WL[338] BL BLB SRAM
    X339 VDD GND WL[339] BL BLB SRAM
    X340 VDD GND WL[340] BL BLB SRAM
    X341 VDD GND WL[341] BL BLB SRAM
    X342 VDD GND WL[342] BL BLB SRAM
    X343 VDD GND WL[343] BL BLB SRAM
    X344 VDD GND WL[344] BL BLB SRAM
    X345 VDD GND WL[345] BL BLB SRAM
    X346 VDD GND WL[346] BL BLB SRAM
    X347 VDD GND WL[347] BL BLB SRAM
    X348 VDD GND WL[348] BL BLB SRAM
    X349 VDD GND WL[349] BL BLB SRAM
    X350 VDD GND WL[350] BL BLB SRAM
    X351 VDD GND WL[351] BL BLB SRAM
    X352 VDD GND WL[352] BL BLB SRAM
    X353 VDD GND WL[353] BL BLB SRAM
    X354 VDD GND WL[354] BL BLB SRAM
    X355 VDD GND WL[355] BL BLB SRAM
    X356 VDD GND WL[356] BL BLB SRAM
    X357 VDD GND WL[357] BL BLB SRAM
    X358 VDD GND WL[358] BL BLB SRAM
    X359 VDD GND WL[359] BL BLB SRAM
    X360 VDD GND WL[360] BL BLB SRAM
    X361 VDD GND WL[361] BL BLB SRAM
    X362 VDD GND WL[362] BL BLB SRAM
    X363 VDD GND WL[363] BL BLB SRAM
    X364 VDD GND WL[364] BL BLB SRAM
    X365 VDD GND WL[365] BL BLB SRAM
    X366 VDD GND WL[366] BL BLB SRAM
    X367 VDD GND WL[367] BL BLB SRAM
    X368 VDD GND WL[368] BL BLB SRAM
    X369 VDD GND WL[369] BL BLB SRAM
    X370 VDD GND WL[370] BL BLB SRAM
    X371 VDD GND WL[371] BL BLB SRAM
    X372 VDD GND WL[372] BL BLB SRAM
    X373 VDD GND WL[373] BL BLB SRAM
    X374 VDD GND WL[374] BL BLB SRAM
    X375 VDD GND WL[375] BL BLB SRAM
    X376 VDD GND WL[376] BL BLB SRAM
    X377 VDD GND WL[377] BL BLB SRAM
    X378 VDD GND WL[378] BL BLB SRAM
    X379 VDD GND WL[379] BL BLB SRAM
    X380 VDD GND WL[380] BL BLB SRAM
    X381 VDD GND WL[381] BL BLB SRAM
    X382 VDD GND WL[382] BL BLB SRAM
    X383 VDD GND WL[383] BL BLB SRAM
    X384 VDD GND WL[384] BL BLB SRAM
    X385 VDD GND WL[385] BL BLB SRAM
    X386 VDD GND WL[386] BL BLB SRAM
    X387 VDD GND WL[387] BL BLB SRAM
    X388 VDD GND WL[388] BL BLB SRAM
    X389 VDD GND WL[389] BL BLB SRAM
    X390 VDD GND WL[390] BL BLB SRAM
    X391 VDD GND WL[391] BL BLB SRAM
    X392 VDD GND WL[392] BL BLB SRAM
    X393 VDD GND WL[393] BL BLB SRAM
    X394 VDD GND WL[394] BL BLB SRAM
    X395 VDD GND WL[395] BL BLB SRAM
    X396 VDD GND WL[396] BL BLB SRAM
    X397 VDD GND WL[397] BL BLB SRAM
    X398 VDD GND WL[398] BL BLB SRAM
    X399 VDD GND WL[399] BL BLB SRAM
    X400 VDD GND WL[400] BL BLB SRAM
    X401 VDD GND WL[401] BL BLB SRAM
    X402 VDD GND WL[402] BL BLB SRAM
    X403 VDD GND WL[403] BL BLB SRAM
    X404 VDD GND WL[404] BL BLB SRAM
    X405 VDD GND WL[405] BL BLB SRAM
    X406 VDD GND WL[406] BL BLB SRAM
    X407 VDD GND WL[407] BL BLB SRAM
    X408 VDD GND WL[408] BL BLB SRAM
    X409 VDD GND WL[409] BL BLB SRAM
    X410 VDD GND WL[410] BL BLB SRAM
    X411 VDD GND WL[411] BL BLB SRAM
    X412 VDD GND WL[412] BL BLB SRAM
    X413 VDD GND WL[413] BL BLB SRAM
    X414 VDD GND WL[414] BL BLB SRAM
    X415 VDD GND WL[415] BL BLB SRAM
    X416 VDD GND WL[416] BL BLB SRAM
    X417 VDD GND WL[417] BL BLB SRAM
    X418 VDD GND WL[418] BL BLB SRAM
    X419 VDD GND WL[419] BL BLB SRAM
    X420 VDD GND WL[420] BL BLB SRAM
    X421 VDD GND WL[421] BL BLB SRAM
    X422 VDD GND WL[422] BL BLB SRAM
    X423 VDD GND WL[423] BL BLB SRAM
    X424 VDD GND WL[424] BL BLB SRAM
    X425 VDD GND WL[425] BL BLB SRAM
    X426 VDD GND WL[426] BL BLB SRAM
    X427 VDD GND WL[427] BL BLB SRAM
    X428 VDD GND WL[428] BL BLB SRAM
    X429 VDD GND WL[429] BL BLB SRAM
    X430 VDD GND WL[430] BL BLB SRAM
    X431 VDD GND WL[431] BL BLB SRAM
    X432 VDD GND WL[432] BL BLB SRAM
    X433 VDD GND WL[433] BL BLB SRAM
    X434 VDD GND WL[434] BL BLB SRAM
    X435 VDD GND WL[435] BL BLB SRAM
    X436 VDD GND WL[436] BL BLB SRAM
    X437 VDD GND WL[437] BL BLB SRAM
    X438 VDD GND WL[438] BL BLB SRAM
    X439 VDD GND WL[439] BL BLB SRAM
    X440 VDD GND WL[440] BL BLB SRAM
    X441 VDD GND WL[441] BL BLB SRAM
    X442 VDD GND WL[442] BL BLB SRAM
    X443 VDD GND WL[443] BL BLB SRAM
    X444 VDD GND WL[444] BL BLB SRAM
    X445 VDD GND WL[445] BL BLB SRAM
    X446 VDD GND WL[446] BL BLB SRAM
    X447 VDD GND WL[447] BL BLB SRAM
    X448 VDD GND WL[448] BL BLB SRAM
    X449 VDD GND WL[449] BL BLB SRAM
    X450 VDD GND WL[450] BL BLB SRAM
    X451 VDD GND WL[451] BL BLB SRAM
    X452 VDD GND WL[452] BL BLB SRAM
    X453 VDD GND WL[453] BL BLB SRAM
    X454 VDD GND WL[454] BL BLB SRAM
    X455 VDD GND WL[455] BL BLB SRAM
    X456 VDD GND WL[456] BL BLB SRAM
    X457 VDD GND WL[457] BL BLB SRAM
    X458 VDD GND WL[458] BL BLB SRAM
    X459 VDD GND WL[459] BL BLB SRAM
    X460 VDD GND WL[460] BL BLB SRAM
    X461 VDD GND WL[461] BL BLB SRAM
    X462 VDD GND WL[462] BL BLB SRAM
    X463 VDD GND WL[463] BL BLB SRAM
    X464 VDD GND WL[464] BL BLB SRAM
    X465 VDD GND WL[465] BL BLB SRAM
    X466 VDD GND WL[466] BL BLB SRAM
    X467 VDD GND WL[467] BL BLB SRAM
    X468 VDD GND WL[468] BL BLB SRAM
    X469 VDD GND WL[469] BL BLB SRAM
    X470 VDD GND WL[470] BL BLB SRAM
    X471 VDD GND WL[471] BL BLB SRAM
    X472 VDD GND WL[472] BL BLB SRAM
    X473 VDD GND WL[473] BL BLB SRAM
    X474 VDD GND WL[474] BL BLB SRAM
    X475 VDD GND WL[475] BL BLB SRAM
    X476 VDD GND WL[476] BL BLB SRAM
    X477 VDD GND WL[477] BL BLB SRAM
    X478 VDD GND WL[478] BL BLB SRAM
    X479 VDD GND WL[479] BL BLB SRAM
    X480 VDD GND WL[480] BL BLB SRAM
    X481 VDD GND WL[481] BL BLB SRAM
    X482 VDD GND WL[482] BL BLB SRAM
    X483 VDD GND WL[483] BL BLB SRAM
    X484 VDD GND WL[484] BL BLB SRAM
    X485 VDD GND WL[485] BL BLB SRAM
    X486 VDD GND WL[486] BL BLB SRAM
    X487 VDD GND WL[487] BL BLB SRAM
    X488 VDD GND WL[488] BL BLB SRAM
    X489 VDD GND WL[489] BL BLB SRAM
    X490 VDD GND WL[490] BL BLB SRAM
    X491 VDD GND WL[491] BL BLB SRAM
    X492 VDD GND WL[492] BL BLB SRAM
    X493 VDD GND WL[493] BL BLB SRAM
    X494 VDD GND WL[494] BL BLB SRAM
    X495 VDD GND WL[495] BL BLB SRAM
    X496 VDD GND WL[496] BL BLB SRAM
    X497 VDD GND WL[497] BL BLB SRAM
    X498 VDD GND WL[498] BL BLB SRAM
    X499 VDD GND WL[499] BL BLB SRAM
    X500 VDD GND WL[500] BL BLB SRAM
    X501 VDD GND WL[501] BL BLB SRAM
    X502 VDD GND WL[502] BL BLB SRAM
    X503 VDD GND WL[503] BL BLB SRAM
    X504 VDD GND WL[504] BL BLB SRAM
    X505 VDD GND WL[505] BL BLB SRAM
    X506 VDD GND WL[506] BL BLB SRAM
    X507 VDD GND WL[507] BL BLB SRAM
    X508 VDD GND WL[508] BL BLB SRAM
    X509 VDD GND WL[509] BL BLB SRAM
    X510 VDD GND WL[510] BL BLB SRAM
    X511 VDD GND WL[511] BL BLB SRAM
XSA SEN BL BLB dout doutb SA
CL0  BL GND load
CL1 BLB GND load
*****************************
**     Voltage Source      **
*****************************
.global VDD GND 
.param supply = 0.7v
VVDD VDD GND supply
VCSEL C_SEL GND supply
//load
.PARAM  load = 80f
//clock for 1GHz wuth 50% duty cycle and 0.05ns rise and fall time
Vclk CLK GND PULSE(0 supply 0.45n 0.05n 0.05n 0.5n 1n)
//precharge signal
Vpre PRE GND PULSE(0 supply 0.45n 0.05n 0.05n 0.5n 1n)
//SEN signal
Vsen SEN GND PULSE(0 supply 0.75n 0.05n 0.05n 0.25n 1n)
//WL voltage
VWL0 WL[0] GND PULSE(0 supply 0.45n 0.05n 0.05n 0.5n 1n)
//WL1-WL511
    VWL1 WL[1] GND 0
    VWL2 WL[2] GND 0
    VWL3 WL[3] GND 0
    VWL4 WL[4] GND 0
    VWL5 WL[5] GND 0
    VWL6 WL[6] GND 0
    VWL7 WL[7] GND 0
    VWL8 WL[8] GND 0
    VWL9 WL[9] GND 0
    VWL10 WL[10] GND 0
    VWL11 WL[11] GND 0
    VWL12 WL[12] GND 0
    VWL13 WL[13] GND 0
    VWL14 WL[14] GND 0
    VWL15 WL[15] GND 0
    VWL16 WL[16] GND 0
    VWL17 WL[17] GND 0
    VWL18 WL[18] GND 0
    VWL19 WL[19] GND 0
    VWL20 WL[20] GND 0
    VWL21 WL[21] GND 0
    VWL22 WL[22] GND 0
    VWL23 WL[23] GND 0
    VWL24 WL[24] GND 0
    VWL25 WL[25] GND 0
    VWL26 WL[26] GND 0
    VWL27 WL[27] GND 0
    VWL28 WL[28] GND 0
    VWL29 WL[29] GND 0
    VWL30 WL[30] GND 0
    VWL31 WL[31] GND 0
    VWL32 WL[32] GND 0
    VWL33 WL[33] GND 0
    VWL34 WL[34] GND 0
    VWL35 WL[35] GND 0
    VWL36 WL[36] GND 0
    VWL37 WL[37] GND 0
    VWL38 WL[38] GND 0
    VWL39 WL[39] GND 0
    VWL40 WL[40] GND 0
    VWL41 WL[41] GND 0
    VWL42 WL[42] GND 0
    VWL43 WL[43] GND 0
    VWL44 WL[44] GND 0
    VWL45 WL[45] GND 0
    VWL46 WL[46] GND 0
    VWL47 WL[47] GND 0
    VWL48 WL[48] GND 0
    VWL49 WL[49] GND 0
    VWL50 WL[50] GND 0
    VWL51 WL[51] GND 0
    VWL52 WL[52] GND 0
    VWL53 WL[53] GND 0
    VWL54 WL[54] GND 0
    VWL55 WL[55] GND 0
    VWL56 WL[56] GND 0
    VWL57 WL[57] GND 0
    VWL58 WL[58] GND 0
    VWL59 WL[59] GND 0
    VWL60 WL[60] GND 0
    VWL61 WL[61] GND 0
    VWL62 WL[62] GND 0
    VWL63 WL[63] GND 0
    VWL64 WL[64] GND 0
    VWL65 WL[65] GND 0
    VWL66 WL[66] GND 0
    VWL67 WL[67] GND 0
    VWL68 WL[68] GND 0
    VWL69 WL[69] GND 0
    VWL70 WL[70] GND 0
    VWL71 WL[71] GND 0
    VWL72 WL[72] GND 0
    VWL73 WL[73] GND 0
    VWL74 WL[74] GND 0
    VWL75 WL[75] GND 0
    VWL76 WL[76] GND 0
    VWL77 WL[77] GND 0
    VWL78 WL[78] GND 0
    VWL79 WL[79] GND 0
    VWL80 WL[80] GND 0
    VWL81 WL[81] GND 0
    VWL82 WL[82] GND 0
    VWL83 WL[83] GND 0
    VWL84 WL[84] GND 0
    VWL85 WL[85] GND 0
    VWL86 WL[86] GND 0
    VWL87 WL[87] GND 0
    VWL88 WL[88] GND 0
    VWL89 WL[89] GND 0
    VWL90 WL[90] GND 0
    VWL91 WL[91] GND 0
    VWL92 WL[92] GND 0
    VWL93 WL[93] GND 0
    VWL94 WL[94] GND 0
    VWL95 WL[95] GND 0
    VWL96 WL[96] GND 0
    VWL97 WL[97] GND 0
    VWL98 WL[98] GND 0
    VWL99 WL[99] GND 0
    VWL100 WL[100] GND 0
    VWL101 WL[101] GND 0
    VWL102 WL[102] GND 0
    VWL103 WL[103] GND 0
    VWL104 WL[104] GND 0
    VWL105 WL[105] GND 0
    VWL106 WL[106] GND 0
    VWL107 WL[107] GND 0
    VWL108 WL[108] GND 0
    VWL109 WL[109] GND 0
    VWL110 WL[110] GND 0
    VWL111 WL[111] GND 0
    VWL112 WL[112] GND 0
    VWL113 WL[113] GND 0
    VWL114 WL[114] GND 0
    VWL115 WL[115] GND 0
    VWL116 WL[116] GND 0
    VWL117 WL[117] GND 0
    VWL118 WL[118] GND 0
    VWL119 WL[119] GND 0
    VWL120 WL[120] GND 0
    VWL121 WL[121] GND 0
    VWL122 WL[122] GND 0
    VWL123 WL[123] GND 0
    VWL124 WL[124] GND 0
    VWL125 WL[125] GND 0
    VWL126 WL[126] GND 0
    VWL127 WL[127] GND 0
    VWL128 WL[128] GND 0
    VWL129 WL[129] GND 0
    VWL130 WL[130] GND 0
    VWL131 WL[131] GND 0
    VWL132 WL[132] GND 0
    VWL133 WL[133] GND 0
    VWL134 WL[134] GND 0
    VWL135 WL[135] GND 0
    VWL136 WL[136] GND 0
    VWL137 WL[137] GND 0
    VWL138 WL[138] GND 0
    VWL139 WL[139] GND 0
    VWL140 WL[140] GND 0
    VWL141 WL[141] GND 0
    VWL142 WL[142] GND 0
    VWL143 WL[143] GND 0
    VWL144 WL[144] GND 0
    VWL145 WL[145] GND 0
    VWL146 WL[146] GND 0
    VWL147 WL[147] GND 0
    VWL148 WL[148] GND 0
    VWL149 WL[149] GND 0
    VWL150 WL[150] GND 0
    VWL151 WL[151] GND 0
    VWL152 WL[152] GND 0
    VWL153 WL[153] GND 0
    VWL154 WL[154] GND 0
    VWL155 WL[155] GND 0
    VWL156 WL[156] GND 0
    VWL157 WL[157] GND 0
    VWL158 WL[158] GND 0
    VWL159 WL[159] GND 0
    VWL160 WL[160] GND 0
    VWL161 WL[161] GND 0
    VWL162 WL[162] GND 0
    VWL163 WL[163] GND 0
    VWL164 WL[164] GND 0
    VWL165 WL[165] GND 0
    VWL166 WL[166] GND 0
    VWL167 WL[167] GND 0
    VWL168 WL[168] GND 0
    VWL169 WL[169] GND 0
    VWL170 WL[170] GND 0
    VWL171 WL[171] GND 0
    VWL172 WL[172] GND 0
    VWL173 WL[173] GND 0
    VWL174 WL[174] GND 0
    VWL175 WL[175] GND 0
    VWL176 WL[176] GND 0
    VWL177 WL[177] GND 0
    VWL178 WL[178] GND 0
    VWL179 WL[179] GND 0
    VWL180 WL[180] GND 0
    VWL181 WL[181] GND 0
    VWL182 WL[182] GND 0
    VWL183 WL[183] GND 0
    VWL184 WL[184] GND 0
    VWL185 WL[185] GND 0
    VWL186 WL[186] GND 0
    VWL187 WL[187] GND 0
    VWL188 WL[188] GND 0
    VWL189 WL[189] GND 0
    VWL190 WL[190] GND 0
    VWL191 WL[191] GND 0
    VWL192 WL[192] GND 0
    VWL193 WL[193] GND 0
    VWL194 WL[194] GND 0
    VWL195 WL[195] GND 0
    VWL196 WL[196] GND 0
    VWL197 WL[197] GND 0
    VWL198 WL[198] GND 0
    VWL199 WL[199] GND 0
    VWL200 WL[200] GND 0
    VWL201 WL[201] GND 0
    VWL202 WL[202] GND 0
    VWL203 WL[203] GND 0
    VWL204 WL[204] GND 0
    VWL205 WL[205] GND 0
    VWL206 WL[206] GND 0
    VWL207 WL[207] GND 0
    VWL208 WL[208] GND 0
    VWL209 WL[209] GND 0
    VWL210 WL[210] GND 0
    VWL211 WL[211] GND 0
    VWL212 WL[212] GND 0
    VWL213 WL[213] GND 0
    VWL214 WL[214] GND 0
    VWL215 WL[215] GND 0
    VWL216 WL[216] GND 0
    VWL217 WL[217] GND 0
    VWL218 WL[218] GND 0
    VWL219 WL[219] GND 0
    VWL220 WL[220] GND 0
    VWL221 WL[221] GND 0
    VWL222 WL[222] GND 0
    VWL223 WL[223] GND 0
    VWL224 WL[224] GND 0
    VWL225 WL[225] GND 0
    VWL226 WL[226] GND 0
    VWL227 WL[227] GND 0
    VWL228 WL[228] GND 0
    VWL229 WL[229] GND 0
    VWL230 WL[230] GND 0
    VWL231 WL[231] GND 0
    VWL232 WL[232] GND 0
    VWL233 WL[233] GND 0
    VWL234 WL[234] GND 0
    VWL235 WL[235] GND 0
    VWL236 WL[236] GND 0
    VWL237 WL[237] GND 0
    VWL238 WL[238] GND 0
    VWL239 WL[239] GND 0
    VWL240 WL[240] GND 0
    VWL241 WL[241] GND 0
    VWL242 WL[242] GND 0
    VWL243 WL[243] GND 0
    VWL244 WL[244] GND 0
    VWL245 WL[245] GND 0
    VWL246 WL[246] GND 0
    VWL247 WL[247] GND 0
    VWL248 WL[248] GND 0
    VWL249 WL[249] GND 0
    VWL250 WL[250] GND 0
    VWL251 WL[251] GND 0
    VWL252 WL[252] GND 0
    VWL253 WL[253] GND 0
    VWL254 WL[254] GND 0
    VWL255 WL[255] GND 0
    VWL256 WL[256] GND 0
    VWL257 WL[257] GND 0
    VWL258 WL[258] GND 0
    VWL259 WL[259] GND 0
    VWL260 WL[260] GND 0
    VWL261 WL[261] GND 0
    VWL262 WL[262] GND 0
    VWL263 WL[263] GND 0
    VWL264 WL[264] GND 0
    VWL265 WL[265] GND 0
    VWL266 WL[266] GND 0
    VWL267 WL[267] GND 0
    VWL268 WL[268] GND 0
    VWL269 WL[269] GND 0
    VWL270 WL[270] GND 0
    VWL271 WL[271] GND 0
    VWL272 WL[272] GND 0
    VWL273 WL[273] GND 0
    VWL274 WL[274] GND 0
    VWL275 WL[275] GND 0
    VWL276 WL[276] GND 0
    VWL277 WL[277] GND 0
    VWL278 WL[278] GND 0
    VWL279 WL[279] GND 0
    VWL280 WL[280] GND 0
    VWL281 WL[281] GND 0
    VWL282 WL[282] GND 0
    VWL283 WL[283] GND 0
    VWL284 WL[284] GND 0
    VWL285 WL[285] GND 0
    VWL286 WL[286] GND 0
    VWL287 WL[287] GND 0
    VWL288 WL[288] GND 0
    VWL289 WL[289] GND 0
    VWL290 WL[290] GND 0
    VWL291 WL[291] GND 0
    VWL292 WL[292] GND 0
    VWL293 WL[293] GND 0
    VWL294 WL[294] GND 0
    VWL295 WL[295] GND 0
    VWL296 WL[296] GND 0
    VWL297 WL[297] GND 0
    VWL298 WL[298] GND 0
    VWL299 WL[299] GND 0
    VWL300 WL[300] GND 0
    VWL301 WL[301] GND 0
    VWL302 WL[302] GND 0
    VWL303 WL[303] GND 0
    VWL304 WL[304] GND 0
    VWL305 WL[305] GND 0
    VWL306 WL[306] GND 0
    VWL307 WL[307] GND 0
    VWL308 WL[308] GND 0
    VWL309 WL[309] GND 0
    VWL310 WL[310] GND 0
    VWL311 WL[311] GND 0
    VWL312 WL[312] GND 0
    VWL313 WL[313] GND 0
    VWL314 WL[314] GND 0
    VWL315 WL[315] GND 0
    VWL316 WL[316] GND 0
    VWL317 WL[317] GND 0
    VWL318 WL[318] GND 0
    VWL319 WL[319] GND 0
    VWL320 WL[320] GND 0
    VWL321 WL[321] GND 0
    VWL322 WL[322] GND 0
    VWL323 WL[323] GND 0
    VWL324 WL[324] GND 0
    VWL325 WL[325] GND 0
    VWL326 WL[326] GND 0
    VWL327 WL[327] GND 0
    VWL328 WL[328] GND 0
    VWL329 WL[329] GND 0
    VWL330 WL[330] GND 0
    VWL331 WL[331] GND 0
    VWL332 WL[332] GND 0
    VWL333 WL[333] GND 0
    VWL334 WL[334] GND 0
    VWL335 WL[335] GND 0
    VWL336 WL[336] GND 0
    VWL337 WL[337] GND 0
    VWL338 WL[338] GND 0
    VWL339 WL[339] GND 0
    VWL340 WL[340] GND 0
    VWL341 WL[341] GND 0
    VWL342 WL[342] GND 0
    VWL343 WL[343] GND 0
    VWL344 WL[344] GND 0
    VWL345 WL[345] GND 0
    VWL346 WL[346] GND 0
    VWL347 WL[347] GND 0
    VWL348 WL[348] GND 0
    VWL349 WL[349] GND 0
    VWL350 WL[350] GND 0
    VWL351 WL[351] GND 0
    VWL352 WL[352] GND 0
    VWL353 WL[353] GND 0
    VWL354 WL[354] GND 0
    VWL355 WL[355] GND 0
    VWL356 WL[356] GND 0
    VWL357 WL[357] GND 0
    VWL358 WL[358] GND 0
    VWL359 WL[359] GND 0
    VWL360 WL[360] GND 0
    VWL361 WL[361] GND 0
    VWL362 WL[362] GND 0
    VWL363 WL[363] GND 0
    VWL364 WL[364] GND 0
    VWL365 WL[365] GND 0
    VWL366 WL[366] GND 0
    VWL367 WL[367] GND 0
    VWL368 WL[368] GND 0
    VWL369 WL[369] GND 0
    VWL370 WL[370] GND 0
    VWL371 WL[371] GND 0
    VWL372 WL[372] GND 0
    VWL373 WL[373] GND 0
    VWL374 WL[374] GND 0
    VWL375 WL[375] GND 0
    VWL376 WL[376] GND 0
    VWL377 WL[377] GND 0
    VWL378 WL[378] GND 0
    VWL379 WL[379] GND 0
    VWL380 WL[380] GND 0
    VWL381 WL[381] GND 0
    VWL382 WL[382] GND 0
    VWL383 WL[383] GND 0
    VWL384 WL[384] GND 0
    VWL385 WL[385] GND 0
    VWL386 WL[386] GND 0
    VWL387 WL[387] GND 0
    VWL388 WL[388] GND 0
    VWL389 WL[389] GND 0
    VWL390 WL[390] GND 0
    VWL391 WL[391] GND 0
    VWL392 WL[392] GND 0
    VWL393 WL[393] GND 0
    VWL394 WL[394] GND 0
    VWL395 WL[395] GND 0
    VWL396 WL[396] GND 0
    VWL397 WL[397] GND 0
    VWL398 WL[398] GND 0
    VWL399 WL[399] GND 0
    VWL400 WL[400] GND 0
    VWL401 WL[401] GND 0
    VWL402 WL[402] GND 0
    VWL403 WL[403] GND 0
    VWL404 WL[404] GND 0
    VWL405 WL[405] GND 0
    VWL406 WL[406] GND 0
    VWL407 WL[407] GND 0
    VWL408 WL[408] GND 0
    VWL409 WL[409] GND 0
    VWL410 WL[410] GND 0
    VWL411 WL[411] GND 0
    VWL412 WL[412] GND 0
    VWL413 WL[413] GND 0
    VWL414 WL[414] GND 0
    VWL415 WL[415] GND 0
    VWL416 WL[416] GND 0
    VWL417 WL[417] GND 0
    VWL418 WL[418] GND 0
    VWL419 WL[419] GND 0
    VWL420 WL[420] GND 0
    VWL421 WL[421] GND 0
    VWL422 WL[422] GND 0
    VWL423 WL[423] GND 0
    VWL424 WL[424] GND 0
    VWL425 WL[425] GND 0
    VWL426 WL[426] GND 0
    VWL427 WL[427] GND 0
    VWL428 WL[428] GND 0
    VWL429 WL[429] GND 0
    VWL430 WL[430] GND 0
    VWL431 WL[431] GND 0
    VWL432 WL[432] GND 0
    VWL433 WL[433] GND 0
    VWL434 WL[434] GND 0
    VWL435 WL[435] GND 0
    VWL436 WL[436] GND 0
    VWL437 WL[437] GND 0
    VWL438 WL[438] GND 0
    VWL439 WL[439] GND 0
    VWL440 WL[440] GND 0
    VWL441 WL[441] GND 0
    VWL442 WL[442] GND 0
    VWL443 WL[443] GND 0
    VWL444 WL[444] GND 0
    VWL445 WL[445] GND 0
    VWL446 WL[446] GND 0
    VWL447 WL[447] GND 0
    VWL448 WL[448] GND 0
    VWL449 WL[449] GND 0
    VWL450 WL[450] GND 0
    VWL451 WL[451] GND 0
    VWL452 WL[452] GND 0
    VWL453 WL[453] GND 0
    VWL454 WL[454] GND 0
    VWL455 WL[455] GND 0
    VWL456 WL[456] GND 0
    VWL457 WL[457] GND 0
    VWL458 WL[458] GND 0
    VWL459 WL[459] GND 0
    VWL460 WL[460] GND 0
    VWL461 WL[461] GND 0
    VWL462 WL[462] GND 0
    VWL463 WL[463] GND 0
    VWL464 WL[464] GND 0
    VWL465 WL[465] GND 0
    VWL466 WL[466] GND 0
    VWL467 WL[467] GND 0
    VWL468 WL[468] GND 0
    VWL469 WL[469] GND 0
    VWL470 WL[470] GND 0
    VWL471 WL[471] GND 0
    VWL472 WL[472] GND 0
    VWL473 WL[473] GND 0
    VWL474 WL[474] GND 0
    VWL475 WL[475] GND 0
    VWL476 WL[476] GND 0
    VWL477 WL[477] GND 0
    VWL478 WL[478] GND 0
    VWL479 WL[479] GND 0
    VWL480 WL[480] GND 0
    VWL481 WL[481] GND 0
    VWL482 WL[482] GND 0
    VWL483 WL[483] GND 0
    VWL484 WL[484] GND 0
    VWL485 WL[485] GND 0
    VWL486 WL[486] GND 0
    VWL487 WL[487] GND 0
    VWL488 WL[488] GND 0
    VWL489 WL[489] GND 0
    VWL490 WL[490] GND 0
    VWL491 WL[491] GND 0
    VWL492 WL[492] GND 0
    VWL493 WL[493] GND 0
    VWL494 WL[494] GND 0
    VWL495 WL[495] GND 0
    VWL496 WL[496] GND 0
    VWL497 WL[497] GND 0
    VWL498 WL[498] GND 0
    VWL499 WL[499] GND 0
    VWL500 WL[500] GND 0
    VWL501 WL[501] GND 0
    VWL502 WL[502] GND 0
    VWL503 WL[503] GND 0
    VWL504 WL[504] GND 0
    VWL505 WL[505] GND 0
    VWL506 WL[506] GND 0
    VWL507 WL[507] GND 0
    VWL508 WL[508] GND 0
    VWL509 WL[509] GND 0
    VWL510 WL[510] GND 0
    VWL511 WL[511] GND 0

***-----------------------***
***       simulation      *** 
***-----------------------***
    .tran 0.1n 10n
*****************************
**    Simulator setting    **
*****************************
    .option post 
    .options probe
    .op
    .probe v(*) i(*)

    .TEMP 25
*****************************
**      Measurement        ** 
*****************************
//power consumption
.meas tran avg_power avg power from=0.1ns to=10ns 
//read access time
.meas tran read_access_time trig v(WL[0]) val='supply/2' targ v(dout) val='supply/2'
***-----------------------***
***      sub-circuit      ***
***-----------------------***
//6T SRAM cell
.subckt SRAM VDD GND WL BL BLB
    Mpr  q   qb  VDD  x  pmos_sram  m=1
    Mnr  q   qb  GND  x  nmos_sram  m=1

    Mpl  qb  q  VDD  x  pmos_sram  m=1
    Mnl  qb  q  GND  x  nmos_sram  m=1

    Mnpr BL  WL  q    x  nmos_sram  m=1
    Mnpl BLB WL  qb   x  nmos_sram  m=1
.ends
//SA
.subckt SA SEN BL BLB O1 O2
    Mp0 O1 SEN BL  BL  pmos_rvt m=1
    Mp1 O2 SEN BLB BLB pmos_rvt m=1

    Mpl O2 O1 VDD VDD pmos_rvt m=1
    Mnl O2 O1 n0  n0  nmos_rvt m=1

    Mpr O1 O2 VDD VDD pmos_rvt m=1
    Mnr O1 O2 n0  n0  nmos_rvt m=1

    Men n0 SEN GND GND nmos_rvt m=1
.ends
.end
